`ifndef SHA256TYPES_VH
    `define SHA256TYPES_VH
    `define WORD [31:0]
    `define LONG [63:0]
`endif